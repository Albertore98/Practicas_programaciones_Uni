library IEEE;
use IEEE.std